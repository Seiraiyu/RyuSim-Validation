// IEEE 1800-2023 Section 11.4.7 - Logical operators
module logical (
    input  logic [7:0] a, b,
    output logic       and_out, or_out, not_out
);
    assign and_out = a && b;
    assign or_out  = a || b;
    assign not_out = !a;
endmodule
