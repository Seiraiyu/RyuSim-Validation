// IEEE 1800-2023 Section 9.4.2 - Sequential logic with asynchronous reset
module d_ff_async_rst (
    input  logic clk,
    input  logic rst_n,
    input  logic d,
    output logic q
);
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            q <= 1'b0;
        else
            q <= d;
    end
endmodule
